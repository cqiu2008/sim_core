////////////////////////////////////////////////////////////////////////////////////////////////////
//  
//  TASKS 
//  
////////////////////////////////////////////////////////////////////////////////////////////////////

////////////////////////////////////////////////////////////////////////////////////////////////////
//  reset 
////////////////////////////////////////////////////////////////////////////////////////////////////
task reset;
  begin

  end
endtask

