`timescale 1ns / 1ps
//`define IPEN  1

//`define ALLCRU 
  `define PERICRU 

module tb_dut_top;
////////////////////////////////////////////////////////////////////////////////////////////////////
//  Common  
////////////////////////////////////////////////////////////////////////////////////////////////////
reg[1024*8:1] msg = 0               ;

always @( msg ) begin
  //$display("[%t] %0s",$realtime,msg);
  $display("\033[1;45m [%t] %0s \033[0m",$realtime,msg);
end
////////////////////////////////////////////////////////////////////////////////////////////////////
//  Environment 
////////////////////////////////////////////////////////////////////////////////////////////////////
`ifdef ALLCRU
  `include "cru/envcru.vh"
`endif
`ifdef PERICRU
  `include "cru_peri/envcru_peri.vh"
`endif

////////////////////////////////////////////////////////////////////////////////////////////////////
//  Tasks
////////////////////////////////////////////////////////////////////////////////////////////////////
// task clkdly(bit [31:0]num, ref logic inter_clk);
//   begin
//     repeat(num)begin
//       @(posedge inter_clk);
//     end
//     #1;
//   end
// endtask

`ifdef ALLCRU
  `include "cru/tskcru.vh"
`endif
`ifdef PERICRU
  `include "cru_peri/tskcru_peri.vh"
`endif

////////////////////////////////////////////////////////////////////////////////////////////////////
//  Testcase 
////////////////////////////////////////////////////////////////////////////////////////////////////
`ifdef ALLCRU
  `include "cru/tccru.vh"
`endif
`ifdef PERICRU 
  `include "cru_peri/tccru_peri.vh"
`endif

////////////////////////////////////////////////////////////////////////////////////////////////////
//  generate fsdb	
////////////////////////////////////////////////////////////////////////////////////////////////////
initial begin
  $fsdbDumpvars("+fsdbfile+tb_dut_top.fsdb");
	$fsdbDumpMDA;
  $fsdbDumpSVA;
end

endmodule

