package e1_pkg;

	import uvm_pkg::*;
	`include "uvm_macros.svh"
	`include "utb/config/e1_config.sv"
	`include "utb/agent/e1_agent/e1_seq_item.sv"
	`include "utb/agent/e1_agent/e1_input_monitor.sv"
	`include "utb/agent/e1_agent/e1_output_monitor.sv"
	`include "utb/agent/e1_agent/e1_input_sequencer.sv"
	`include "utb/agent/e1_agent/e1_input_seq.sv"
	`include "utb/agent/e1_agent/e1_input_driver.sv"
	`include "utb/agent/e1_agent/e1_agent.sv"


endpackage
