////////////////////////////////////////////////////////////////////////////////////////////////////
//  xxx testcase  
////////////////////////////////////////////////////////////////////////////////////////////////////
integer i;

initial begin

  //This test creates four errors
  //force tb_dut_top.uut.uut_0.ERR_MAX_INT = 4;
  
  #55;  
  //reset 
  //reset;
  //standby(100);
end
