//--------------------------------------------------------------------------------------------------
//File Name    : rclk_and_rrst_tsk 
//Author       : qiu.chao 
//--------------------------------------------------------------------------------------------------
//Module Hierarchy :
//rclk_and_rrst_tsk_inst |-rclk_and_rrst_tsk
//--------------------------------------------------------------------------------------------------
//Release History :
//Version         Date           Author        Description
// 1.0          2019-01-01       qiu.chao       1st draft
//--------------------------------------------------------------------------------------------------
//Main Function Tree:
//a)rclk_and_rrst_tsk: 
//Description Function:
//rclk_and_rrst_tsk
//--------------------------------------------------------------------------------------------------

////////////////////////////////////////////////////////////////////////////////////////////////////
// Naming specification																			  // 
////////////////////////////////////////////////////////////////////////////////////////////////////

////////////////////////////////////////////////////////////////////////////////////////////////////
//		rclk generator
////////////////////////////////////////////////////////////////////////////////////////////////////
initial begin
	rclk = 0;
end
always #19 rclk =~rclk;

////////////////////////////////////////////////////////////////////////////////////////////////////
//		rrst task
////////////////////////////////////////////////////////////////////////////////////////////////////
initial begin
	rrst = 0; 
end

task rrst_tsk;
input [31:0]rst_num;
begin
	rrst = 1'b0;
	repeat (1) @(posedge rclk);
	#1
	rrst = 1'b1;
	repeat (rst_num) @(posedge rclk);
	#1
	rrst = 1'b0;
	repeat (1) @(posedge rclk);
	#1;
end
endtask

////////////////////////////////////////////////////////////////////////////////////////////////////
//                                                                                                //
//    __    __    __    __    __    __    __    __    __    __    __    __    __    __    __    __//
// __|  |__|  |__|  |__|  |__|  |__|  |__|  |__|  |__|  |__|  |__|  |__|  |__|  |__|  |__|  |__|  |/
//                                                                                                //
//                                                                                                //
////////////////////////////////////////////////////////////////////////////////////////////////////
