package eth_pkg;

	import uvm_pkg::*;
	`include "uvm_macros.svh"
	`include "utb/config/eth_public_config.sv"
	`include "utb/config/eth_private_config.sv"
	`include "utb/agent/eth_agent/eth_seq_item.sv"
	`include "utb/agent/eth_agent/eth_output_monitor.sv"
	`include "utb/agent/eth_agent/eth_input_sequencer.sv"
	`include "utb/agent/eth_agent/eth_input_seq.sv"
	`include "utb/agent/eth_agent/eth_input_driver.sv"
	`include "utb/agent/eth_agent/eth_agent.sv"

endpackage
