//--------------------------------------------------------------------------------------------------
//File Name    : xxx 
//Author       : xxx 
//--------------------------------------------------------------------------------------------------
//Module Hierarchy :
//xxx_inst |-xxx
//--------------------------------------------------------------------------------------------------
//Release History :
//Version         Date           Author        Description
// 1.0          2019-01-01       xxx			1st draft
//--------------------------------------------------------------------------------------------------
//Main Function Tree:
//a)xxx: 
//Description Function:
//xxx
//--------------------------------------------------------------------------------------------------
module xxx();
////////////////////////////////////////////////////////////////////////////////////////////////////
// Naming specification																			  // 
// (1)																							  // 
////////////////////////////////////////////////////////////////////////////////////////////////////

////////////////////////////////////////////////////////////////////////////////////////////////////
//                                                                                                //
//    __    __    __    __    __    __    __    __    __    __    __    __    __    __    __    __//
// __|  |__|  |__|  |__|  |__|  |__|  |__|  |__|  |__|  |__|  |__|  |__|  |__|  |__|  |__|  |__|  |/
//                                                                                                //
//                                                                                                //
////////////////////////////////////////////////////////////////////////////////////////////////////

////////////////////////////////////////////////////////////////////////////////////////////////////
//		xxx_name																				  //	
////////////////////////////////////////////////////////////////////////////////////////////////////

endmodule

