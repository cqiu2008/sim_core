`timescale 1ns / 1ps
//`define IPEN  1

module tb_dut_top;
////////////////////////////////////////////////////////////////////////////////////////////////////
//  Common  
////////////////////////////////////////////////////////////////////////////////////////////////////
reg         npor                          ;// i                    
reg         soc_test_mode                 ;// i
reg         soc_scan_mode                 ;// i
reg         soc_mbist_mode                ;// i
reg         scan_clk_ahb                  ;// i
reg         scan_clk_apb                  ;// i
reg         scan_clk_func                 ;// i
reg         chiprstn_top                  ;// i

initial begin
  npor            <= 0 ;// i                    
  soc_test_mode   <= 0 ;// i
  soc_scan_mode   <= 0 ;// i
  soc_mbist_mode  <= 0 ;// i
  scan_clk_ahb    <= 0 ;// i
  scan_clk_apb    <= 0 ;// i
  scan_clk_func   <= 0 ;// i
  chiprstn_top    <= 0 ;// i
end

////////////////////////////////////////////////////////////////////////////////////////////////////
//  Environment 
////////////////////////////////////////////////////////////////////////////////////////////////////
`include "envcru_peri.vh"

////////////////////////////////////////////////////////////////////////////////////////////////////
//  Tasks
////////////////////////////////////////////////////////////////////////////////////////////////////
`include "tskcru_peri.vh"

////////////////////////////////////////////////////////////////////////////////////////////////////
//  Testcase 
////////////////////////////////////////////////////////////////////////////////////////////////////
`include "tccru_peri.vh"

////////////////////////////////////////////////////////////////////////////////////////////////////
//  generate fsdb	
////////////////////////////////////////////////////////////////////////////////////////////////////
initial begin
  $fsdbDumpvars("+fsdbfile+tb_dut_top.fsdb");
	$fsdbDumpMDA;
  $fsdbDumpSVA;
end

endmodule

